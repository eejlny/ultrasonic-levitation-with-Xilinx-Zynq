library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_UltrasonicLogic is
generic(
    Trans : integer := 64
    );
end tb_UltrasonicLogic;

architecture Behavioral of tb_UltrasonicLogic is

component UltrasonicLogic is
  generic(
    TRANSDUCER_NUM : integer := 64
    );
  Port (   
           Emmitter_clk : in STD_LOGIC; 
           Control : in STD_LOGIC_VECTOR(3 downto 0);
           Match : in STD_LOGIC_VECTOR ((8*Trans)-1 downto 0);
           Mask : in std_logic_vector(Trans-1 downto 0);
           Phases : out STD_LOGIC_VECTOR (Trans-1 downto 0);
           Sync : out std_logic
           );
end component UltrasonicLogic;

signal tb_MATCH: STD_LOGIC_VECTOR((8*Trans)-1 downto 0);

signal tb_RST : STD_LOGIC := '1';
signal tb_CHANNEL_VALUES: STD_LOGIC_VECTOR(Trans-1 downto 0);
signal tb_CTRL : std_logic_vector(3 downto 0);
signal tb_sync : std_logic;
signal tb_leds : std_logic_vector(1 downto 0);

signal tb_AXI_CLK : std_logic := '0';
signal tb_CLK : STD_LOGIC := '0';

signal tb_Mask :std_logic_vector(Trans-1 downto 0) := "0000000000000000000000000000000011111111111111111111111111111111";



begin
tb_CLK <= not tb_CLK after 48828.125 ps;
tb_AXI_CLK <= not tb_AXI_CLK after 5000 ps;
tb_RST <= '1';



mapping:UltrasonicLogic
generic map(
    TRANSDUCER_NUM => Trans
    )
port map(
    
    Emmitter_clk => tb_CLK,
    Control => tb_CTRL,
    Match => tb_MATCH, 
    Phases => tb_CHANNEL_VALUES,
    Mask => tb_Mask,
    Sync => tb_sync
);

process
begin
tb_MATCH <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

wait for 781250 ps;
tb_CTRL <= "0000";
wait for 781250 ps;
tb_CTRL <= "1111";
wait for 100 us;
tb_MATCH <= "00000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000000";
wait for 100 us;
tb_MATCH <= "11111111111111101111110111111100111110111111101011111001111110001111011111110110111101011111010011110011111100101111000111110000111011111110111011101101111011001110101111101010111010011110100011100111111001101110010111100100111000111110001011100001111000001101111111011110110111011101110011011011110110101101100111011000110101111101011011010101110101001101001111010010110100011101000011001111110011101100110111001100110010111100101011001001110010001100011111000110110001011100010011000011110000101100000111000000";
wait for 100 us;
tb_CTRL <= "0000";
wait for 100 us;
tb_CTRL <= "0001";
wait for 100 us;
tb_CTRL <= "0010";
wait for 100 us;
tb_CTRL <= "0011";
wait for 100 us;
tb_CTRL <= "0100";
wait for 100 us;
tb_CTRL <= "0101";
wait for 100 us;
tb_CTRL <= "0110";
wait for 100 us;
tb_CTRL <= "0111";
wait for 100 us;
tb_CTRL <= "1000";
wait for 100 us;
tb_CTRL <= "1001";
wait for 100 us;
tb_CTRL <= "1010";
wait for 100 us;
tb_CTRL <= "1011";
wait for 100 us;
tb_CTRL <= "1100";
wait for 100 us;
tb_CTRL <= "1101";
wait for 100 us;
tb_CTRL <= "1110";
wait for 100 us;
tb_CTRL <= "1111";



--tb_MATCH <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--wait for 100 us;
--tb_MATCH <= "0010111101001011110000101110110010111010001011100100101110000010110111001011011000101101010010110100001011001100101100100010110001001011000000101011110010101110001010110100101011000010101011001010101000101010010010101000001010011100101001100010100101001010010000101000110010100010001010000100101000000010011111001001111000100111010010011100001001101100100110100010011001001001100000100101110010010110001001010100100101000010010011001001001000100100010010010000001000111100100011100010001101001000110000100010110010001010001000100100100010000010000111001000011000100001010010000100001000001100100000100010000001001000000000011111110001111110";
--wait for 100 us;
--tb_MATCH <= "0011111100001111101100111110100011111001001111100000111101110011110110001111010100111101000011110011001111001000111100010011110000001110111100111011100011101101001110110000111010110011101010001110100100111010000011100111001110011000111001010011100100001110001100111000100011100001001110000000110111110011011110001101110100110111000011011011001101101000110110010011011000001101011100110101100011010101001101010000110100110011010010001101000100110100000011001111001100111000110011010011001100001100101100110010100011001001001100100000110001110011000110001100010100110001000011000011001100001000110000010011000000001011111100101111100010111101";
--wait for 100 us;
--tb_MATCH <= "0100111011010011101001001110010100111000010011011101001101100100110101010011010001001100110100110010010011000101001100000100101111010010111001001011010100101100010010101101001010100100101001010010100001001001110100100110010010010101001001000100100011010010001001001000010100100000010001111101000111100100011101010001110001000110110100011010010001100101000110000100010111010001011001000101010100010100010001001101000100100100010001010001000001000011110100001110010000110101000011000100001011010000101001000010010100001000010000011101000001100100000101010000010001000000110100000010010000000101000000000011111111001111111000111111010011111100";
--wait for 100 us;
--tb_MATCH <= "0101111010010111100101011110000101110111010111011001011101010101110100010111001101011100100101110001010111000001011011110101101110010110110101011011000101101011010110101001011010010101101000010110011101011001100101100101010110010001011000110101100010010110000101011000000101011111010101111001010111010101011100010101101101010110100101011001010101100001010101110101010110010101010101010101000101010011010101001001010100010101010000010100111101010011100101001101010100110001010010110101001010010100100101010010000101000111010100011001010001010101000100010100001101010000100101000001010100000001001111110100111110010011110101001111000100111011";
--wait for 100 us;
--tb_MATCH <= "0110111001011011100001101101110110110110011011010101101101000110110011011011001001101100010110110000011010111101101011100110101101011010110001101010110110101010011010100101101010000110100111011010011001101001010110100100011010001101101000100110100001011010000001100111110110011110011001110101100111000110011011011001101001100110010110011000011001011101100101100110010101011001010001100100110110010010011001000101100100000110001111011000111001100011010110001100011000101101100010100110001001011000100001100001110110000110011000010101100001000110000011011000001001100000010110000000010111111101011111100101111101010111110001011110110101111010";
--wait for 100 us;
--tb_MATCH <= "0111111000011111011101111101100111110101011111010001111100110111110010011111000101111100000111101111011110111001111011010111101100011110101101111010100111101001011110100001111001110111100110011110010101111001000111100011011110001001111000010111100000011101111101110111100111011101011101110001110110110111011010011101100101110110000111010111011101011001110101010111010100011101001101110100100111010001011101000001110011110111001110011100110101110011000111001011011100101001110010010111001000011100011101110001100111000101011100010001110000110111000010011100000101110000000110111111011011111001101111010110111100011011101101101110100110111001";
--wait for 100 us;
--tb_MATCH <= "1000110111100011011010001101011000110100100011001110001100101000110001100011000010001011111000101110100010110110001011001000101011100010101010001010011000101000100010011110001001101000100101100010010010001000111000100010100010000110001000001000011111100001111010000111011000011100100001101110000110101000011001100001100010000101111000010110100001010110000101001000010011100001001010000100011000010000100000111110000011101000001101100000110010000010111000001010100000100110000010001000000111100000011010000001011000000100100000001110000000101000000001100000000001111111110111111110011111110101111111000111111011011111101001111110010111111000";
--wait for 100 us;
--tb_MATCH <= "1001110110100111010110011101001001110011100111001010011100011001110000100110111110011011101001101101100110110010011010111001101010100110100110011010001001100111100110011010011001011001100100100110001110011000101001100001100110000010010111111001011110100101110110010111001001011011100101101010010110011001011000100101011110010101101001010101100101010010010100111001010010100101000110010100001001001111100100111010010011011001001100100100101110010010101001001001100100100010010001111001000110100100010110010001001001000011100100001010010000011001000000100011111110001111101000111101100011110010001110111000111010100011100110001110001000110111";
--wait for 100 us;
--tb_MATCH <= "1010110101101011010010101100111010110010101011000110101100001010101111101010111010101011011010101100101010101110101010101010101001101010100010101001111010100110101010010110101001001010100011101010001010101000011010100000101001111110100111101010011101101001110010100110111010011010101001100110100110001010010111101001011010100101011010010100101001001110100100101010010001101001000010100011111010001110101000110110100011001010001011101000101010100010011010001000101000011110100001101010000101101000010010100000111010000010101000000110100000001001111111100111111010011111011001111100100111101110011110101001111001100111100010011101111001110110";
--wait for 100 us;
--tb_MATCH <= "1011110100101111001110111100101011110001101111000010111011111011101110101110110110111011001011101011101110101010111010011011101000101110011110111001101011100101101110010010111000111011100010101110000110111000001011011111101101111010110111011011011100101101101110110110101011011001101101100010110101111011010110101101010110110101001011010011101101001010110100011011010000101100111110110011101011001101101100110010110010111011001010101100100110110010001011000111101100011010110001011011000100101100001110110000101011000001101100000010101111111010111110101011110110101111001010111011101011101010101110011010111000101011011110101101101010110101";
--wait for 100 us;
--tb_MATCH <= "1100110011110011001011001100011100110000110010111111001011101100101101110010110011001010111100101010110010100111001010001100100111110010011011001001011100100100110010001111001000101100100001110010000011000111111100011110110001110111000111001100011011110001101011000110011100011000110001011111000101101100010101110001010011000100111100010010110001000111000100001100001111110000111011000011011100001100110000101111000010101100001001110000100011000001111100000110110000010111000001001100000011110000001011000000011100000000101111111110111111101011111101101111110010111110111011111010101111100110111110001011110111101111011010111101011011110100";
--wait for 100 us;
--tb_MATCH <= "1101110010110111000111011100001101101111110110111011011011011101101100110110101111011010101101101001110110100011011001111101100110110110010111011001001101100011110110001011011000011101100000110101111111010111101101011101110101110011010110111101011010110101100111010110001101010111110101011011010101011101010100110101001111010100101101010001110101000011010011111101001110110100110111010011001101001011110100101011010010011101001000110100011111010001101101000101110100010011010000111101000010110100000111010000001100111111110011111011001111011100111100110011101111001110101100111001110011100011001101111100110110110011010111001101001100110011";
--wait for 100 us;
--tb_MATCH <= "1110110010111011000111101100001110101111111010111011101011011110101100111010101111101010101110101001111010100011101001111110100110111010010111101001001110100011111010001011101000011110100000111001111111100111101110011101111001110011100110111110011010111001100111100110001110010111111001011011100101011110010100111001001111100100101110010001111001000011100011111110001110111000110111100011001110001011111000101011100010011110001000111000011111100001101110000101111000010011100000111110000010111000000111100000001101111111110111111011011111011101111100110111101111011110101101111001110111100011011101111101110110110111010111011101001101110011";
--wait for 100 us;
--tb_MATCH <= "1111110001111111000011111011111111101110111110110111111011001111101011111110101011111010011111101000111110011111111001101111100101111110010011111000111111100010111110000111111000001111011111111101111011110111011111011100111101101111110110101111011001111101100011110101111111010110111101010111110101001111010011111101001011110100011111010000111100111111110011101111001101111100110011110010111111001010111100100111110010001111000111111100011011110001011111000100111100001111110000101111000001111100000011101111111110111110111011110111101111001110111011111011101011101110011110111000111011011111101101101110110101111011010011101100111110110010";
--wait for 100 us;
--tb_MATCH <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111101111111110011111110111111111010111111100111111110001111110111111111011011111101011111110100111111001111111100101111110001";
--wait for 100 us;
--tb_MATCH <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--wait for 100 us;






loop
wait for 1 ns;
end loop;

end process;


end Behavioral;
